magic
tech sky130A
magscale 1 2
timestamp 1756228627
<< error_p >>
rect -845 181 -787 187
rect -653 181 -595 187
rect -461 181 -403 187
rect -269 181 -211 187
rect -77 181 -19 187
rect 115 181 173 187
rect 307 181 365 187
rect 499 181 557 187
rect 691 181 749 187
rect 883 181 941 187
rect -845 147 -833 181
rect -653 147 -641 181
rect -461 147 -449 181
rect -269 147 -257 181
rect -77 147 -65 181
rect 115 147 127 181
rect 307 147 319 181
rect 499 147 511 181
rect 691 147 703 181
rect 883 147 895 181
rect -845 141 -787 147
rect -653 141 -595 147
rect -461 141 -403 147
rect -269 141 -211 147
rect -77 141 -19 147
rect 115 141 173 147
rect 307 141 365 147
rect 499 141 557 147
rect 691 141 749 147
rect 883 141 941 147
rect -941 -147 -883 -141
rect -749 -147 -691 -141
rect -557 -147 -499 -141
rect -365 -147 -307 -141
rect -173 -147 -115 -141
rect 19 -147 77 -141
rect 211 -147 269 -141
rect 403 -147 461 -141
rect 595 -147 653 -141
rect 787 -147 845 -141
rect -941 -181 -929 -147
rect -749 -181 -737 -147
rect -557 -181 -545 -147
rect -365 -181 -353 -147
rect -173 -181 -161 -147
rect 19 -181 31 -147
rect 211 -181 223 -147
rect 403 -181 415 -147
rect 595 -181 607 -147
rect 787 -181 799 -147
rect -941 -187 -883 -181
rect -749 -187 -691 -181
rect -557 -187 -499 -181
rect -365 -187 -307 -181
rect -173 -187 -115 -181
rect 19 -187 77 -181
rect 211 -187 269 -181
rect 403 -187 461 -181
rect 595 -187 653 -181
rect 787 -187 845 -181
<< nwell >>
rect -1127 -319 1127 319
<< pmos >>
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
<< pdiff >>
rect -989 88 -927 100
rect -989 -88 -977 88
rect -943 -88 -927 88
rect -989 -100 -927 -88
rect -897 88 -831 100
rect -897 -88 -881 88
rect -847 -88 -831 88
rect -897 -100 -831 -88
rect -801 88 -735 100
rect -801 -88 -785 88
rect -751 -88 -735 88
rect -801 -100 -735 -88
rect -705 88 -639 100
rect -705 -88 -689 88
rect -655 -88 -639 88
rect -705 -100 -639 -88
rect -609 88 -543 100
rect -609 -88 -593 88
rect -559 -88 -543 88
rect -609 -100 -543 -88
rect -513 88 -447 100
rect -513 -88 -497 88
rect -463 -88 -447 88
rect -513 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 513 100
rect 447 -88 463 88
rect 497 -88 513 88
rect 447 -100 513 -88
rect 543 88 609 100
rect 543 -88 559 88
rect 593 -88 609 88
rect 543 -100 609 -88
rect 639 88 705 100
rect 639 -88 655 88
rect 689 -88 705 88
rect 639 -100 705 -88
rect 735 88 801 100
rect 735 -88 751 88
rect 785 -88 801 88
rect 735 -100 801 -88
rect 831 88 897 100
rect 831 -88 847 88
rect 881 -88 897 88
rect 831 -100 897 -88
rect 927 88 989 100
rect 927 -88 943 88
rect 977 -88 989 88
rect 927 -100 989 -88
<< pdiffc >>
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
<< nsubdiff >>
rect -1091 249 -995 283
rect 995 249 1091 283
rect -1091 187 -1057 249
rect 1057 187 1091 249
rect -1091 -249 -1057 -187
rect 1057 -249 1091 -187
rect -1091 -283 -995 -249
rect 995 -283 1091 -249
<< nsubdiffcont >>
rect -995 249 995 283
rect -1091 -187 -1057 187
rect 1057 -187 1091 187
rect -995 -283 995 -249
<< poly >>
rect -849 181 -783 197
rect -849 147 -833 181
rect -799 147 -783 181
rect -849 131 -783 147
rect -657 181 -591 197
rect -657 147 -641 181
rect -607 147 -591 181
rect -657 131 -591 147
rect -465 181 -399 197
rect -465 147 -449 181
rect -415 147 -399 181
rect -465 131 -399 147
rect -273 181 -207 197
rect -273 147 -257 181
rect -223 147 -207 181
rect -273 131 -207 147
rect -81 181 -15 197
rect -81 147 -65 181
rect -31 147 -15 181
rect -81 131 -15 147
rect 111 181 177 197
rect 111 147 127 181
rect 161 147 177 181
rect 111 131 177 147
rect 303 181 369 197
rect 303 147 319 181
rect 353 147 369 181
rect 303 131 369 147
rect 495 181 561 197
rect 495 147 511 181
rect 545 147 561 181
rect 495 131 561 147
rect 687 181 753 197
rect 687 147 703 181
rect 737 147 753 181
rect 687 131 753 147
rect 879 181 945 197
rect 879 147 895 181
rect 929 147 945 181
rect 879 131 945 147
rect -927 100 -897 126
rect -831 100 -801 131
rect -735 100 -705 126
rect -639 100 -609 131
rect -543 100 -513 126
rect -447 100 -417 131
rect -351 100 -321 126
rect -255 100 -225 131
rect -159 100 -129 126
rect -63 100 -33 131
rect 33 100 63 126
rect 129 100 159 131
rect 225 100 255 126
rect 321 100 351 131
rect 417 100 447 126
rect 513 100 543 131
rect 609 100 639 126
rect 705 100 735 131
rect 801 100 831 126
rect 897 100 927 131
rect -927 -131 -897 -100
rect -831 -126 -801 -100
rect -735 -131 -705 -100
rect -639 -126 -609 -100
rect -543 -131 -513 -100
rect -447 -126 -417 -100
rect -351 -131 -321 -100
rect -255 -126 -225 -100
rect -159 -131 -129 -100
rect -63 -126 -33 -100
rect 33 -131 63 -100
rect 129 -126 159 -100
rect 225 -131 255 -100
rect 321 -126 351 -100
rect 417 -131 447 -100
rect 513 -126 543 -100
rect 609 -131 639 -100
rect 705 -126 735 -100
rect 801 -131 831 -100
rect 897 -126 927 -100
rect -945 -147 -879 -131
rect -945 -181 -929 -147
rect -895 -181 -879 -147
rect -945 -197 -879 -181
rect -753 -147 -687 -131
rect -753 -181 -737 -147
rect -703 -181 -687 -147
rect -753 -197 -687 -181
rect -561 -147 -495 -131
rect -561 -181 -545 -147
rect -511 -181 -495 -147
rect -561 -197 -495 -181
rect -369 -147 -303 -131
rect -369 -181 -353 -147
rect -319 -181 -303 -147
rect -369 -197 -303 -181
rect -177 -147 -111 -131
rect -177 -181 -161 -147
rect -127 -181 -111 -147
rect -177 -197 -111 -181
rect 15 -147 81 -131
rect 15 -181 31 -147
rect 65 -181 81 -147
rect 15 -197 81 -181
rect 207 -147 273 -131
rect 207 -181 223 -147
rect 257 -181 273 -147
rect 207 -197 273 -181
rect 399 -147 465 -131
rect 399 -181 415 -147
rect 449 -181 465 -147
rect 399 -197 465 -181
rect 591 -147 657 -131
rect 591 -181 607 -147
rect 641 -181 657 -147
rect 591 -197 657 -181
rect 783 -147 849 -131
rect 783 -181 799 -147
rect 833 -181 849 -147
rect 783 -197 849 -181
<< polycont >>
rect -833 147 -799 181
rect -641 147 -607 181
rect -449 147 -415 181
rect -257 147 -223 181
rect -65 147 -31 181
rect 127 147 161 181
rect 319 147 353 181
rect 511 147 545 181
rect 703 147 737 181
rect 895 147 929 181
rect -929 -181 -895 -147
rect -737 -181 -703 -147
rect -545 -181 -511 -147
rect -353 -181 -319 -147
rect -161 -181 -127 -147
rect 31 -181 65 -147
rect 223 -181 257 -147
rect 415 -181 449 -147
rect 607 -181 641 -147
rect 799 -181 833 -147
<< locali >>
rect -1091 249 -995 283
rect 995 249 1091 283
rect -1091 187 -1057 249
rect 1057 187 1091 249
rect -849 147 -833 181
rect -799 147 -783 181
rect -657 147 -641 181
rect -607 147 -591 181
rect -465 147 -449 181
rect -415 147 -399 181
rect -273 147 -257 181
rect -223 147 -207 181
rect -81 147 -65 181
rect -31 147 -15 181
rect 111 147 127 181
rect 161 147 177 181
rect 303 147 319 181
rect 353 147 369 181
rect 495 147 511 181
rect 545 147 561 181
rect 687 147 703 181
rect 737 147 753 181
rect 879 147 895 181
rect 929 147 945 181
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -881 88 -847 104
rect -881 -104 -847 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -689 88 -655 104
rect -689 -104 -655 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 655 88 689 104
rect 655 -104 689 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 847 88 881 104
rect 847 -104 881 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect -945 -181 -929 -147
rect -895 -181 -879 -147
rect -753 -181 -737 -147
rect -703 -181 -687 -147
rect -561 -181 -545 -147
rect -511 -181 -495 -147
rect -369 -181 -353 -147
rect -319 -181 -303 -147
rect -177 -181 -161 -147
rect -127 -181 -111 -147
rect 15 -181 31 -147
rect 65 -181 81 -147
rect 207 -181 223 -147
rect 257 -181 273 -147
rect 399 -181 415 -147
rect 449 -181 465 -147
rect 591 -181 607 -147
rect 641 -181 657 -147
rect 783 -181 799 -147
rect 833 -181 849 -147
rect -1091 -249 -1057 -187
rect 1057 -249 1091 -187
rect -1091 -283 -995 -249
rect 995 -283 1091 -249
<< viali >>
rect -833 147 -799 181
rect -641 147 -607 181
rect -449 147 -415 181
rect -257 147 -223 181
rect -65 147 -31 181
rect 127 147 161 181
rect 319 147 353 181
rect 511 147 545 181
rect 703 147 737 181
rect 895 147 929 181
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect -929 -181 -895 -147
rect -737 -181 -703 -147
rect -545 -181 -511 -147
rect -353 -181 -319 -147
rect -161 -181 -127 -147
rect 31 -181 65 -147
rect 223 -181 257 -147
rect 415 -181 449 -147
rect 607 -181 641 -147
rect 799 -181 833 -147
<< metal1 >>
rect -845 181 -787 187
rect -845 147 -833 181
rect -799 147 -787 181
rect -845 141 -787 147
rect -653 181 -595 187
rect -653 147 -641 181
rect -607 147 -595 181
rect -653 141 -595 147
rect -461 181 -403 187
rect -461 147 -449 181
rect -415 147 -403 181
rect -461 141 -403 147
rect -269 181 -211 187
rect -269 147 -257 181
rect -223 147 -211 181
rect -269 141 -211 147
rect -77 181 -19 187
rect -77 147 -65 181
rect -31 147 -19 181
rect -77 141 -19 147
rect 115 181 173 187
rect 115 147 127 181
rect 161 147 173 181
rect 115 141 173 147
rect 307 181 365 187
rect 307 147 319 181
rect 353 147 365 181
rect 307 141 365 147
rect 499 181 557 187
rect 499 147 511 181
rect 545 147 557 181
rect 499 141 557 147
rect 691 181 749 187
rect 691 147 703 181
rect 737 147 749 181
rect 691 141 749 147
rect 883 181 941 187
rect 883 147 895 181
rect 929 147 941 181
rect 883 141 941 147
rect -983 88 -937 100
rect -983 -88 -977 88
rect -943 -88 -937 88
rect -983 -100 -937 -88
rect -887 88 -841 100
rect -887 -88 -881 88
rect -847 -88 -841 88
rect -887 -100 -841 -88
rect -791 88 -745 100
rect -791 -88 -785 88
rect -751 -88 -745 88
rect -791 -100 -745 -88
rect -695 88 -649 100
rect -695 -88 -689 88
rect -655 -88 -649 88
rect -695 -100 -649 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 649 88 695 100
rect 649 -88 655 88
rect 689 -88 695 88
rect 649 -100 695 -88
rect 745 88 791 100
rect 745 -88 751 88
rect 785 -88 791 88
rect 745 -100 791 -88
rect 841 88 887 100
rect 841 -88 847 88
rect 881 -88 887 88
rect 841 -100 887 -88
rect 937 88 983 100
rect 937 -88 943 88
rect 977 -88 983 88
rect 937 -100 983 -88
rect -941 -147 -883 -141
rect -941 -181 -929 -147
rect -895 -181 -883 -147
rect -941 -187 -883 -181
rect -749 -147 -691 -141
rect -749 -181 -737 -147
rect -703 -181 -691 -147
rect -749 -187 -691 -181
rect -557 -147 -499 -141
rect -557 -181 -545 -147
rect -511 -181 -499 -147
rect -557 -187 -499 -181
rect -365 -147 -307 -141
rect -365 -181 -353 -147
rect -319 -181 -307 -147
rect -365 -187 -307 -181
rect -173 -147 -115 -141
rect -173 -181 -161 -147
rect -127 -181 -115 -147
rect -173 -187 -115 -181
rect 19 -147 77 -141
rect 19 -181 31 -147
rect 65 -181 77 -147
rect 19 -187 77 -181
rect 211 -147 269 -141
rect 211 -181 223 -147
rect 257 -181 269 -147
rect 211 -187 269 -181
rect 403 -147 461 -141
rect 403 -181 415 -147
rect 449 -181 461 -147
rect 403 -187 461 -181
rect 595 -147 653 -141
rect 595 -181 607 -147
rect 641 -181 653 -147
rect 595 -187 653 -181
rect 787 -147 845 -141
rect 787 -181 799 -147
rect 833 -181 845 -147
rect 787 -187 845 -181
<< properties >>
string FIXED_BBOX -1074 -266 1074 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
