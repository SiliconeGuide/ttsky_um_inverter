magic
tech sky130A
magscale 1 2
timestamp 1756927211
<< metal1 >>
rect 10915 6170 11305 6176
rect 11305 5780 22484 6170
rect 10915 5774 11305 5780
rect 20830 4480 22062 4660
rect 26600 4654 26824 4692
rect 20830 4100 21010 4480
rect 26600 4474 27414 4654
rect 26600 4450 26824 4474
rect 26622 4436 26802 4450
rect 20824 3920 20830 4100
rect 21010 3920 21016 4100
rect 27234 3368 27414 4474
rect 21693 3021 22488 3358
rect 27228 3188 27234 3368
rect 27414 3188 27420 3368
rect 18473 2631 18479 3021
rect 18869 2968 22488 3021
rect 18869 2631 22083 2968
<< via1 >>
rect 10915 5780 11305 6170
rect 20830 3920 21010 4100
rect 27234 3188 27414 3368
rect 18479 2631 18869 3021
<< metal2 >>
rect 9322 5780 9331 6170
rect 9721 5780 10915 6170
rect 11305 5780 11311 6170
rect 20830 4100 21010 4106
rect 20830 3397 21010 3920
rect 20830 3227 20835 3397
rect 21005 3227 21010 3397
rect 20830 3222 21010 3227
rect 27234 3368 27414 3374
rect 20835 3218 21005 3222
rect 18479 3021 18869 3027
rect 17560 2631 17569 3021
rect 17959 2631 18479 3021
rect 27234 2697 27414 3188
rect 18479 2625 18869 2631
rect 27230 2527 27239 2697
rect 27409 2527 27418 2697
rect 27234 2522 27414 2527
<< via2 >>
rect 9331 5780 9721 6170
rect 20835 3227 21005 3397
rect 17569 2631 17959 3021
rect 27239 2527 27409 2697
<< metal3 >>
rect 9326 6170 9726 6175
rect 6909 5780 6915 6170
rect 7305 5780 9331 6170
rect 9721 5780 9726 6170
rect 9326 5775 9726 5780
rect 20830 3397 21010 3402
rect 20830 3227 20835 3397
rect 21005 3227 21010 3397
rect 17564 3021 17964 3026
rect 16533 2631 16539 3021
rect 16929 2631 17569 3021
rect 17959 2631 17964 3021
rect 17564 2626 17964 2631
rect 20830 1572 21010 3227
rect 27234 2697 27414 2702
rect 27234 2527 27239 2697
rect 27409 2527 27414 2697
rect 27234 2111 27414 2527
rect 27229 1933 27235 2111
rect 27413 1933 27419 2111
rect 27234 1932 27414 1933
rect 20830 1566 23054 1572
rect 20830 1392 23550 1566
rect 22854 1386 23550 1392
rect 23370 971 23550 1386
rect 23365 793 23371 971
rect 23549 793 23555 971
rect 23370 792 23550 793
<< via3 >>
rect 6915 5780 7305 6170
rect 16539 2631 16929 3021
rect 27235 1933 27413 2111
rect 23371 793 23549 971
<< metal4 >>
rect 3006 44598 3066 45152
rect 3558 44598 3618 45152
rect 4110 44598 4170 45152
rect 4662 44598 4722 45152
rect 5214 44598 5274 45152
rect 5766 44598 5826 45152
rect 6318 44598 6378 45152
rect 6870 44598 6930 45152
rect 7422 44598 7482 45152
rect 7974 44598 8034 45152
rect 8526 44598 8586 45152
rect 9078 44598 9138 45152
rect 9630 44598 9690 45152
rect 10182 44598 10242 45152
rect 10734 44598 10794 45152
rect 11286 44598 11346 45152
rect 11838 44598 11898 45152
rect 12390 44598 12450 45152
rect 12942 44598 13002 45152
rect 13494 44598 13554 45152
rect 14046 44598 14106 45152
rect 14598 44598 14658 45152
rect 15150 44598 15210 45152
rect 15702 44598 15762 45152
rect 16254 44952 16314 45152
rect 16806 44952 16866 45152
rect 17358 44952 17418 45152
rect 17910 44952 17970 45152
rect 18462 44952 18522 45152
rect 19014 44952 19074 45152
rect 19566 44952 19626 45152
rect 20118 44952 20178 45152
rect 20670 44952 20730 45152
rect 21222 44952 21282 45152
rect 21774 44952 21834 45152
rect 22326 44952 22386 45152
rect 22878 44952 22938 45152
rect 23430 44952 23490 45152
rect 23982 44952 24042 45152
rect 24534 44952 24594 45152
rect 25086 44952 25146 45152
rect 25638 44952 25698 45152
rect 26190 44952 26250 45152
rect 244 6170 644 44140
rect 2770 44122 15844 44598
rect 6914 6170 7306 6171
rect 230 5780 6915 6170
rect 7305 5780 7306 6170
rect 244 988 644 5780
rect 6914 5779 7306 5780
rect 13504 3021 13904 44122
rect 16538 3021 16930 3022
rect 13504 2631 16539 3021
rect 16929 2631 16930 3021
rect 13504 1002 13904 2631
rect 16538 2630 16930 2631
rect 27234 2111 27414 2112
rect 27234 1933 27235 2111
rect 27413 1933 27414 2111
rect 23370 971 23550 972
rect 23370 793 23371 971
rect 23549 793 23550 971
rect 186 0 366 200
rect 4050 0 4230 200
rect 7914 0 8094 200
rect 11778 0 11958 200
rect 15642 0 15822 200
rect 19506 0 19686 200
rect 23370 0 23550 793
rect 27234 0 27414 1933
use double_inverter  double_inverter_1
timestamp 1756234663
transform 1 0 21298 0 1 4972
box 492 -2004 5504 1198
<< labels >>
flabel metal4 s 25638 44952 25698 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 26190 44952 26250 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 27234 0 27414 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 23370 0 23550 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 19506 0 19686 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 15642 0 15822 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 11778 0 11958 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 s 7914 0 8094 200 0 FreeSans 960 0 0 0 ua[5]
port 8 nsew signal bidirectional
flabel metal4 s 4050 0 4230 200 0 FreeSans 960 0 0 0 ua[6]
port 9 nsew signal bidirectional
flabel metal4 s 186 0 366 200 0 FreeSans 960 0 0 0 ua[7]
port 10 nsew signal bidirectional
flabel metal4 s 24534 44952 24594 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 11 nsew signal input
flabel metal4 s 23982 44952 24042 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 12 nsew signal input
flabel metal4 s 23430 44952 23490 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 14 nsew signal input
flabel metal4 s 22326 44952 22386 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 15 nsew signal input
flabel metal4 s 21774 44952 21834 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 16 nsew signal input
flabel metal4 s 21222 44952 21282 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 17 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 18 nsew signal input
flabel metal4 s 20118 44952 20178 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 19 nsew signal input
flabel metal4 s 19566 44952 19626 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 20 nsew signal input
flabel metal4 s 19014 44952 19074 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 21 nsew signal input
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 22 nsew signal input
flabel metal4 s 17910 44952 17970 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 23 nsew signal input
flabel metal4 s 17358 44952 17418 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 24 nsew signal input
flabel metal4 s 16806 44952 16866 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 25 nsew signal input
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 26 nsew signal input
flabel metal4 s 6870 44952 6930 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 27 nsew signal output
flabel metal4 s 6318 44952 6378 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 28 nsew signal output
flabel metal4 s 5766 44952 5826 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 29 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 30 nsew signal output
flabel metal4 s 4662 44952 4722 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 31 nsew signal output
flabel metal4 s 4110 44952 4170 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 32 nsew signal output
flabel metal4 s 3558 44952 3618 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 33 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 34 nsew signal output
flabel metal4 s 11286 44952 11346 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 35 nsew signal output
flabel metal4 s 10734 44952 10794 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 36 nsew signal output
flabel metal4 s 10182 44952 10242 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 37 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 38 nsew signal output
flabel metal4 s 9078 44952 9138 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 39 nsew signal output
flabel metal4 s 8526 44952 8586 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 40 nsew signal output
flabel metal4 s 7974 44952 8034 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 41 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 42 nsew signal output
flabel metal4 s 15702 44952 15762 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 43 nsew signal output
flabel metal4 s 15150 44952 15210 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 44 nsew signal output
flabel metal4 s 14598 44952 14658 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 45 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 46 nsew signal output
flabel metal4 s 13494 44952 13554 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 47 nsew signal output
flabel metal4 s 12942 44952 13002 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 48 nsew signal output
flabel metal4 s 12390 44952 12450 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 49 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 50 nsew signal output
flabel metal4 13504 1002 13904 44154 1 FreeSans 1600 0 0 0 VGND
port 52 nsew ground bidirectional
flabel metal4 244 988 644 44140 1 FreeSans 1600 0 0 0 VAPWR
port 53 nsew power bidirectional
<< properties >>
string FIXED_BBOX 0 0 29072 45152
<< end >>
