magic
tech sky130A
magscale 1 2
timestamp 1756182476
<< error_p >>
rect 351 621 386 638
rect 352 620 386 621
rect 352 584 422 620
rect 738 584 791 585
rect 182 553 240 559
rect 182 519 194 553
rect 369 550 440 584
rect 720 550 791 584
rect 182 513 240 519
rect 369 89 439 550
rect 721 549 791 550
rect 738 515 809 549
rect 2921 515 2956 532
rect 551 482 609 488
rect 551 448 563 482
rect 551 442 609 448
rect 551 172 609 178
rect 551 138 563 172
rect 551 132 609 138
rect 369 53 422 89
rect 738 36 808 515
rect 2922 514 2956 515
rect 2922 478 2992 514
rect 1020 447 1078 453
rect 1212 447 1270 453
rect 1404 447 1462 453
rect 1596 447 1654 453
rect 1788 447 1846 453
rect 1980 447 2038 453
rect 2172 447 2230 453
rect 2364 447 2422 453
rect 2556 447 2614 453
rect 2748 447 2806 453
rect 1020 413 1032 447
rect 1212 413 1224 447
rect 1404 413 1416 447
rect 1596 413 1608 447
rect 1788 413 1800 447
rect 1980 413 1992 447
rect 2172 413 2184 447
rect 2364 413 2376 447
rect 2556 413 2568 447
rect 2748 413 2760 447
rect 2939 444 3010 478
rect 1020 407 1078 413
rect 1212 407 1270 413
rect 1404 407 1462 413
rect 1596 407 1654 413
rect 1788 407 1846 413
rect 1980 407 2038 413
rect 2172 407 2230 413
rect 2364 407 2422 413
rect 2556 407 2614 413
rect 2748 407 2806 413
rect 924 119 982 125
rect 1116 119 1174 125
rect 1308 119 1366 125
rect 1500 119 1558 125
rect 1692 119 1750 125
rect 1884 119 1942 125
rect 2076 119 2134 125
rect 2268 119 2326 125
rect 2460 119 2518 125
rect 2652 119 2710 125
rect 924 85 936 119
rect 1116 85 1128 119
rect 1308 85 1320 119
rect 1500 85 1512 119
rect 1692 85 1704 119
rect 1884 85 1896 119
rect 2076 85 2088 119
rect 2268 85 2280 119
rect 2460 85 2472 119
rect 2652 85 2664 119
rect 924 79 982 85
rect 1116 79 1174 85
rect 1308 79 1366 85
rect 1500 79 1558 85
rect 1692 79 1750 85
rect 1884 79 1942 85
rect 2076 79 2134 85
rect 2268 79 2326 85
rect 2460 79 2518 85
rect 2652 79 2710 85
rect 738 0 791 36
rect 2939 -17 3009 444
rect 3221 376 3279 382
rect 3413 376 3471 382
rect 3605 376 3663 382
rect 3797 376 3855 382
rect 3989 376 4047 382
rect 4181 376 4239 382
rect 4373 376 4431 382
rect 4565 376 4623 382
rect 4757 376 4815 382
rect 4949 376 5007 382
rect 3221 342 3233 376
rect 3413 342 3425 376
rect 3605 342 3617 376
rect 3797 342 3809 376
rect 3989 342 4001 376
rect 4181 342 4193 376
rect 4373 342 4385 376
rect 4565 342 4577 376
rect 4757 342 4769 376
rect 4949 342 4961 376
rect 3221 336 3279 342
rect 3413 336 3471 342
rect 3605 336 3663 342
rect 3797 336 3855 342
rect 3989 336 4047 342
rect 4181 336 4239 342
rect 4373 336 4431 342
rect 4565 336 4623 342
rect 4757 336 4815 342
rect 4949 336 5007 342
rect 3125 66 3183 72
rect 3317 66 3375 72
rect 3509 66 3567 72
rect 3701 66 3759 72
rect 3893 66 3951 72
rect 4085 66 4143 72
rect 4277 66 4335 72
rect 4469 66 4527 72
rect 4661 66 4719 72
rect 4853 66 4911 72
rect 3125 32 3137 66
rect 3317 32 3329 66
rect 3509 32 3521 66
rect 3701 32 3713 66
rect 3893 32 3905 66
rect 4085 32 4097 66
rect 4277 32 4289 66
rect 4469 32 4481 66
rect 4661 32 4673 66
rect 4853 32 4865 66
rect 3125 26 3183 32
rect 3317 26 3375 32
rect 3509 26 3567 32
rect 3701 26 3759 32
rect 3893 26 3951 32
rect 4085 26 4143 32
rect 4277 26 4335 32
rect 4469 26 4527 32
rect 4661 26 4719 32
rect 4853 26 4911 32
rect 2939 -53 2992 -17
use double_inverter  x1
timestamp 1756182476
transform 1 0 53 0 1 1412
box -53 -1518 5140 200
<< end >>
