** sch_path: /home/ttuser/projects/ttsky-analog-template/xschem/double_inverter.sch
.subckt double_inverter VDD VSS input output
*.PININFO VDD:B VSS:B input:I output:O
XM1 inverted input VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=1 nf=1 m=1
XM2 inverted input VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM3 output inverted VDD VDD sky130_fd_pr__pfet_01v8 L=0.15 W=20 nf=20 m=1
XM4 output inverted VSS VSS sky130_fd_pr__nfet_01v8 L=0.15 W=20 nf=20 m=1
.ends
.end
