magic
tech sky130A
magscale 1 2
timestamp 1756234663
<< viali >>
rect 2440 484 4414 518
rect 1324 396 1464 432
rect 1340 -1214 1480 -1172
rect 2448 -1270 4420 -1232
<< metal1 >>
rect 796 808 4664 1198
rect 906 264 1004 808
rect 1302 432 1498 808
rect 2422 518 4442 808
rect 4580 634 4664 808
rect 4574 550 4580 634
rect 4664 550 4670 634
rect 2422 484 2440 518
rect 4414 484 4442 518
rect 2422 468 4442 484
rect 1302 396 1324 432
rect 1464 396 1498 432
rect 1302 378 1498 396
rect 1792 412 2008 414
rect 1792 364 4378 412
rect 1792 278 2148 364
rect 906 166 1374 264
rect 1418 158 2148 278
rect 2428 256 2438 316
rect 2490 256 2500 316
rect 2620 256 2630 316
rect 2682 256 2692 316
rect 2812 256 2822 316
rect 2874 256 2884 316
rect 3004 256 3014 316
rect 3066 256 3076 316
rect 3196 256 3206 316
rect 3258 256 3268 316
rect 3388 256 3398 316
rect 3450 256 3460 316
rect 3580 256 3590 316
rect 3642 256 3652 316
rect 3772 256 3782 316
rect 3834 256 3844 316
rect 3964 256 3974 316
rect 4026 256 4036 316
rect 4156 256 4166 316
rect 4218 256 4228 316
rect 4348 256 4358 316
rect 4410 256 4420 316
rect 1792 86 2148 158
rect 2524 136 2534 196
rect 2586 136 2596 196
rect 2716 136 2726 196
rect 2778 136 2788 196
rect 2908 136 2918 196
rect 2970 136 2980 196
rect 3100 136 3110 196
rect 3162 136 3172 196
rect 3292 136 3302 196
rect 3354 136 3364 196
rect 3484 136 3494 196
rect 3546 136 3556 196
rect 3676 136 3686 196
rect 3738 136 3748 196
rect 3868 136 3878 196
rect 3930 136 3940 196
rect 4060 136 4070 196
rect 4122 136 4132 196
rect 4252 136 4262 196
rect 4314 136 4324 196
rect 898 18 1430 74
rect 1792 30 4284 86
rect 898 -306 1098 18
rect 492 -506 1098 -306
rect 898 -792 1098 -506
rect 898 -854 1452 -792
rect 1792 -802 2148 30
rect 5086 -498 5092 -298
rect 5292 -498 5504 -298
rect 1792 -852 4380 -802
rect 1792 -924 2148 -852
rect 900 -1040 1388 -926
rect 900 -1614 1014 -1040
rect 1432 -1044 2148 -924
rect 2436 -946 2446 -886
rect 2498 -946 2508 -886
rect 2628 -946 2638 -886
rect 2690 -946 2700 -886
rect 2820 -946 2830 -886
rect 2882 -946 2892 -886
rect 3012 -946 3022 -886
rect 3074 -946 3084 -886
rect 3204 -946 3214 -886
rect 3266 -946 3276 -886
rect 3396 -946 3406 -886
rect 3458 -946 3468 -886
rect 3588 -946 3598 -886
rect 3650 -946 3660 -886
rect 3780 -946 3790 -886
rect 3842 -946 3852 -886
rect 3972 -946 3982 -886
rect 4034 -946 4044 -886
rect 4164 -946 4174 -886
rect 4226 -946 4236 -886
rect 4356 -946 4366 -886
rect 4418 -946 4428 -886
rect 1792 -1112 2148 -1044
rect 2532 -1076 2542 -1016
rect 2594 -1076 2604 -1016
rect 2724 -1076 2734 -1016
rect 2786 -1076 2796 -1016
rect 2916 -1076 2926 -1016
rect 2978 -1076 2988 -1016
rect 3108 -1076 3118 -1016
rect 3170 -1076 3180 -1016
rect 3300 -1076 3310 -1016
rect 3362 -1076 3372 -1016
rect 3492 -1076 3502 -1016
rect 3554 -1076 3564 -1016
rect 3684 -1076 3694 -1016
rect 3746 -1076 3756 -1016
rect 3876 -1076 3886 -1016
rect 3938 -1076 3948 -1016
rect 4068 -1076 4078 -1016
rect 4130 -1076 4140 -1016
rect 4260 -1076 4270 -1016
rect 4322 -1076 4332 -1016
rect 1320 -1172 1500 -1148
rect 1792 -1160 4286 -1112
rect 1320 -1214 1340 -1172
rect 1480 -1214 1500 -1172
rect 1320 -1614 1500 -1214
rect 2416 -1232 4436 -1218
rect 2416 -1270 2448 -1232
rect 4420 -1270 4436 -1232
rect 2416 -1614 4436 -1270
rect 4694 -1390 4700 -1306
rect 4784 -1390 4790 -1306
rect 4700 -1614 4784 -1390
rect 800 -2004 4784 -1614
<< via1 >>
rect 4580 550 4664 634
rect 2438 256 2490 316
rect 2630 256 2682 316
rect 2822 256 2874 316
rect 3014 256 3066 316
rect 3206 256 3258 316
rect 3398 256 3450 316
rect 3590 256 3642 316
rect 3782 256 3834 316
rect 3974 256 4026 316
rect 4166 256 4218 316
rect 4358 256 4410 316
rect 2534 136 2586 196
rect 2726 136 2778 196
rect 2918 136 2970 196
rect 3110 136 3162 196
rect 3302 136 3354 196
rect 3494 136 3546 196
rect 3686 136 3738 196
rect 3878 136 3930 196
rect 4070 136 4122 196
rect 4262 136 4314 196
rect 5092 -498 5292 -298
rect 2446 -946 2498 -886
rect 2638 -946 2690 -886
rect 2830 -946 2882 -886
rect 3022 -946 3074 -886
rect 3214 -946 3266 -886
rect 3406 -946 3458 -886
rect 3598 -946 3650 -886
rect 3790 -946 3842 -886
rect 3982 -946 4034 -886
rect 4174 -946 4226 -886
rect 4366 -946 4418 -886
rect 2542 -1076 2594 -1016
rect 2734 -1076 2786 -1016
rect 2926 -1076 2978 -1016
rect 3118 -1076 3170 -1016
rect 3310 -1076 3362 -1016
rect 3502 -1076 3554 -1016
rect 3694 -1076 3746 -1016
rect 3886 -1076 3938 -1016
rect 4078 -1076 4130 -1016
rect 4270 -1076 4322 -1016
rect 4700 -1390 4784 -1306
<< metal2 >>
rect 4580 634 4664 640
rect 4580 326 4664 550
rect 2412 316 4664 326
rect 2412 256 2438 316
rect 2490 256 2630 316
rect 2682 256 2822 316
rect 2874 256 3014 316
rect 3066 256 3206 316
rect 3258 256 3398 316
rect 3450 256 3590 316
rect 3642 256 3782 316
rect 3834 256 3974 316
rect 4026 256 4166 316
rect 4218 256 4358 316
rect 4410 256 4664 316
rect 2412 242 4664 256
rect 2508 196 4858 206
rect 2508 136 2534 196
rect 2586 136 2726 196
rect 2778 136 2918 196
rect 2970 136 3110 196
rect 3162 136 3302 196
rect 3354 136 3494 196
rect 3546 136 3686 196
rect 3738 136 3878 196
rect 3930 136 4070 196
rect 4122 136 4262 196
rect 4314 136 4858 196
rect 2508 122 4858 136
rect 4646 -298 4858 122
rect 5092 -298 5292 -292
rect 4646 -498 5092 -298
rect 4646 -876 4858 -498
rect 5092 -504 5292 -498
rect 2420 -886 4858 -876
rect 2420 -946 2446 -886
rect 2498 -946 2638 -886
rect 2690 -946 2830 -886
rect 2882 -946 3022 -886
rect 3074 -946 3214 -886
rect 3266 -946 3406 -886
rect 3458 -946 3598 -886
rect 3650 -946 3790 -886
rect 3842 -946 3982 -886
rect 4034 -946 4174 -886
rect 4226 -946 4366 -886
rect 4418 -946 4858 -886
rect 2420 -960 4858 -946
rect 4658 -962 4858 -960
rect 2516 -1016 4784 -1006
rect 2516 -1076 2542 -1016
rect 2594 -1076 2734 -1016
rect 2786 -1076 2926 -1016
rect 2978 -1076 3118 -1016
rect 3170 -1076 3310 -1016
rect 3362 -1076 3502 -1016
rect 3554 -1076 3694 -1016
rect 3746 -1076 3886 -1016
rect 3938 -1076 4078 -1016
rect 4130 -1076 4270 -1016
rect 4322 -1076 4784 -1016
rect 2516 -1090 4784 -1076
rect 4700 -1306 4784 -1090
rect 4700 -1396 4784 -1390
use sky130_fd_pr__pfet_01v8_8DVCWJ  sky130_fd_pr__pfet_01v8_8DVCWJ_0
timestamp 1756228627
transform 1 0 3425 0 1 223
box -1127 -319 1127 319
use sky130_fd_pr__pfet_01v8_LGS3BL  XM1
timestamp 1756228627
transform 1 0 1397 0 1 176
box -211 -284 211 284
use sky130_fd_pr__nfet_01v8_64Z3AY  XM2
timestamp 1756228627
transform 1 0 1411 0 1 -957
box -211 -279 211 279
use sky130_fd_pr__nfet_01v8_YTLFGX  XM4
timestamp 1756228627
transform 1 0 3433 0 1 -982
box -1127 -310 1127 310
<< labels >>
flabel metal1 900 904 1100 1104 0 FreeSans 256 0 0 0 VDD
port 0 nsew
flabel metal1 898 -1900 1098 -1700 0 FreeSans 256 0 0 0 VSS
port 1 nsew
flabel metal1 492 -506 692 -306 0 FreeSans 256 0 0 0 input
port 2 nsew
flabel metal1 5304 -498 5504 -298 0 FreeSans 256 0 0 0 output
port 3 nsew
<< end >>
