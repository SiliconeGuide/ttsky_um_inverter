magic
tech sky130A
magscale 1 2
timestamp 1756228627
<< error_p >>
rect -845 172 -787 178
rect -653 172 -595 178
rect -461 172 -403 178
rect -269 172 -211 178
rect -77 172 -19 178
rect 115 172 173 178
rect 307 172 365 178
rect 499 172 557 178
rect 691 172 749 178
rect 883 172 941 178
rect -845 138 -833 172
rect -653 138 -641 172
rect -461 138 -449 172
rect -269 138 -257 172
rect -77 138 -65 172
rect 115 138 127 172
rect 307 138 319 172
rect 499 138 511 172
rect 691 138 703 172
rect 883 138 895 172
rect -845 132 -787 138
rect -653 132 -595 138
rect -461 132 -403 138
rect -269 132 -211 138
rect -77 132 -19 138
rect 115 132 173 138
rect 307 132 365 138
rect 499 132 557 138
rect 691 132 749 138
rect 883 132 941 138
rect -941 -138 -883 -132
rect -749 -138 -691 -132
rect -557 -138 -499 -132
rect -365 -138 -307 -132
rect -173 -138 -115 -132
rect 19 -138 77 -132
rect 211 -138 269 -132
rect 403 -138 461 -132
rect 595 -138 653 -132
rect 787 -138 845 -132
rect -941 -172 -929 -138
rect -749 -172 -737 -138
rect -557 -172 -545 -138
rect -365 -172 -353 -138
rect -173 -172 -161 -138
rect 19 -172 31 -138
rect 211 -172 223 -138
rect 403 -172 415 -138
rect 595 -172 607 -138
rect 787 -172 799 -138
rect -941 -178 -883 -172
rect -749 -178 -691 -172
rect -557 -178 -499 -172
rect -365 -178 -307 -172
rect -173 -178 -115 -172
rect 19 -178 77 -172
rect 211 -178 269 -172
rect 403 -178 461 -172
rect 595 -178 653 -172
rect 787 -178 845 -172
<< pwell >>
rect -1127 -310 1127 310
<< nmos >>
rect -927 -100 -897 100
rect -831 -100 -801 100
rect -735 -100 -705 100
rect -639 -100 -609 100
rect -543 -100 -513 100
rect -447 -100 -417 100
rect -351 -100 -321 100
rect -255 -100 -225 100
rect -159 -100 -129 100
rect -63 -100 -33 100
rect 33 -100 63 100
rect 129 -100 159 100
rect 225 -100 255 100
rect 321 -100 351 100
rect 417 -100 447 100
rect 513 -100 543 100
rect 609 -100 639 100
rect 705 -100 735 100
rect 801 -100 831 100
rect 897 -100 927 100
<< ndiff >>
rect -989 88 -927 100
rect -989 -88 -977 88
rect -943 -88 -927 88
rect -989 -100 -927 -88
rect -897 88 -831 100
rect -897 -88 -881 88
rect -847 -88 -831 88
rect -897 -100 -831 -88
rect -801 88 -735 100
rect -801 -88 -785 88
rect -751 -88 -735 88
rect -801 -100 -735 -88
rect -705 88 -639 100
rect -705 -88 -689 88
rect -655 -88 -639 88
rect -705 -100 -639 -88
rect -609 88 -543 100
rect -609 -88 -593 88
rect -559 -88 -543 88
rect -609 -100 -543 -88
rect -513 88 -447 100
rect -513 -88 -497 88
rect -463 -88 -447 88
rect -513 -100 -447 -88
rect -417 88 -351 100
rect -417 -88 -401 88
rect -367 -88 -351 88
rect -417 -100 -351 -88
rect -321 88 -255 100
rect -321 -88 -305 88
rect -271 -88 -255 88
rect -321 -100 -255 -88
rect -225 88 -159 100
rect -225 -88 -209 88
rect -175 -88 -159 88
rect -225 -100 -159 -88
rect -129 88 -63 100
rect -129 -88 -113 88
rect -79 -88 -63 88
rect -129 -100 -63 -88
rect -33 88 33 100
rect -33 -88 -17 88
rect 17 -88 33 88
rect -33 -100 33 -88
rect 63 88 129 100
rect 63 -88 79 88
rect 113 -88 129 88
rect 63 -100 129 -88
rect 159 88 225 100
rect 159 -88 175 88
rect 209 -88 225 88
rect 159 -100 225 -88
rect 255 88 321 100
rect 255 -88 271 88
rect 305 -88 321 88
rect 255 -100 321 -88
rect 351 88 417 100
rect 351 -88 367 88
rect 401 -88 417 88
rect 351 -100 417 -88
rect 447 88 513 100
rect 447 -88 463 88
rect 497 -88 513 88
rect 447 -100 513 -88
rect 543 88 609 100
rect 543 -88 559 88
rect 593 -88 609 88
rect 543 -100 609 -88
rect 639 88 705 100
rect 639 -88 655 88
rect 689 -88 705 88
rect 639 -100 705 -88
rect 735 88 801 100
rect 735 -88 751 88
rect 785 -88 801 88
rect 735 -100 801 -88
rect 831 88 897 100
rect 831 -88 847 88
rect 881 -88 897 88
rect 831 -100 897 -88
rect 927 88 989 100
rect 927 -88 943 88
rect 977 -88 989 88
rect 927 -100 989 -88
<< ndiffc >>
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
<< psubdiff >>
rect -1091 240 -995 274
rect 995 240 1091 274
rect -1091 178 -1057 240
rect 1057 178 1091 240
rect -1091 -240 -1057 -178
rect 1057 -240 1091 -178
rect -1091 -274 -995 -240
rect 995 -274 1091 -240
<< psubdiffcont >>
rect -995 240 995 274
rect -1091 -178 -1057 178
rect 1057 -178 1091 178
rect -995 -274 995 -240
<< poly >>
rect -849 172 -783 188
rect -849 138 -833 172
rect -799 138 -783 172
rect -927 100 -897 126
rect -849 122 -783 138
rect -657 172 -591 188
rect -657 138 -641 172
rect -607 138 -591 172
rect -831 100 -801 122
rect -735 100 -705 126
rect -657 122 -591 138
rect -465 172 -399 188
rect -465 138 -449 172
rect -415 138 -399 172
rect -639 100 -609 122
rect -543 100 -513 126
rect -465 122 -399 138
rect -273 172 -207 188
rect -273 138 -257 172
rect -223 138 -207 172
rect -447 100 -417 122
rect -351 100 -321 126
rect -273 122 -207 138
rect -81 172 -15 188
rect -81 138 -65 172
rect -31 138 -15 172
rect -255 100 -225 122
rect -159 100 -129 126
rect -81 122 -15 138
rect 111 172 177 188
rect 111 138 127 172
rect 161 138 177 172
rect -63 100 -33 122
rect 33 100 63 126
rect 111 122 177 138
rect 303 172 369 188
rect 303 138 319 172
rect 353 138 369 172
rect 129 100 159 122
rect 225 100 255 126
rect 303 122 369 138
rect 495 172 561 188
rect 495 138 511 172
rect 545 138 561 172
rect 321 100 351 122
rect 417 100 447 126
rect 495 122 561 138
rect 687 172 753 188
rect 687 138 703 172
rect 737 138 753 172
rect 513 100 543 122
rect 609 100 639 126
rect 687 122 753 138
rect 879 172 945 188
rect 879 138 895 172
rect 929 138 945 172
rect 705 100 735 122
rect 801 100 831 126
rect 879 122 945 138
rect 897 100 927 122
rect -927 -122 -897 -100
rect -945 -138 -879 -122
rect -831 -126 -801 -100
rect -735 -122 -705 -100
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -945 -188 -879 -172
rect -753 -138 -687 -122
rect -639 -126 -609 -100
rect -543 -122 -513 -100
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -753 -188 -687 -172
rect -561 -138 -495 -122
rect -447 -126 -417 -100
rect -351 -122 -321 -100
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -561 -188 -495 -172
rect -369 -138 -303 -122
rect -255 -126 -225 -100
rect -159 -122 -129 -100
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -369 -188 -303 -172
rect -177 -138 -111 -122
rect -63 -126 -33 -100
rect 33 -122 63 -100
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect -177 -188 -111 -172
rect 15 -138 81 -122
rect 129 -126 159 -100
rect 225 -122 255 -100
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 15 -188 81 -172
rect 207 -138 273 -122
rect 321 -126 351 -100
rect 417 -122 447 -100
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 207 -188 273 -172
rect 399 -138 465 -122
rect 513 -126 543 -100
rect 609 -122 639 -100
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 399 -188 465 -172
rect 591 -138 657 -122
rect 705 -126 735 -100
rect 801 -122 831 -100
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 591 -188 657 -172
rect 783 -138 849 -122
rect 897 -126 927 -100
rect 783 -172 799 -138
rect 833 -172 849 -138
rect 783 -188 849 -172
<< polycont >>
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
<< locali >>
rect -1091 240 -995 274
rect 995 240 1091 274
rect -1091 178 -1057 240
rect 1057 178 1091 240
rect -849 138 -833 172
rect -799 138 -783 172
rect -657 138 -641 172
rect -607 138 -591 172
rect -465 138 -449 172
rect -415 138 -399 172
rect -273 138 -257 172
rect -223 138 -207 172
rect -81 138 -65 172
rect -31 138 -15 172
rect 111 138 127 172
rect 161 138 177 172
rect 303 138 319 172
rect 353 138 369 172
rect 495 138 511 172
rect 545 138 561 172
rect 687 138 703 172
rect 737 138 753 172
rect 879 138 895 172
rect 929 138 945 172
rect -977 88 -943 104
rect -977 -104 -943 -88
rect -881 88 -847 104
rect -881 -104 -847 -88
rect -785 88 -751 104
rect -785 -104 -751 -88
rect -689 88 -655 104
rect -689 -104 -655 -88
rect -593 88 -559 104
rect -593 -104 -559 -88
rect -497 88 -463 104
rect -497 -104 -463 -88
rect -401 88 -367 104
rect -401 -104 -367 -88
rect -305 88 -271 104
rect -305 -104 -271 -88
rect -209 88 -175 104
rect -209 -104 -175 -88
rect -113 88 -79 104
rect -113 -104 -79 -88
rect -17 88 17 104
rect -17 -104 17 -88
rect 79 88 113 104
rect 79 -104 113 -88
rect 175 88 209 104
rect 175 -104 209 -88
rect 271 88 305 104
rect 271 -104 305 -88
rect 367 88 401 104
rect 367 -104 401 -88
rect 463 88 497 104
rect 463 -104 497 -88
rect 559 88 593 104
rect 559 -104 593 -88
rect 655 88 689 104
rect 655 -104 689 -88
rect 751 88 785 104
rect 751 -104 785 -88
rect 847 88 881 104
rect 847 -104 881 -88
rect 943 88 977 104
rect 943 -104 977 -88
rect -945 -172 -929 -138
rect -895 -172 -879 -138
rect -753 -172 -737 -138
rect -703 -172 -687 -138
rect -561 -172 -545 -138
rect -511 -172 -495 -138
rect -369 -172 -353 -138
rect -319 -172 -303 -138
rect -177 -172 -161 -138
rect -127 -172 -111 -138
rect 15 -172 31 -138
rect 65 -172 81 -138
rect 207 -172 223 -138
rect 257 -172 273 -138
rect 399 -172 415 -138
rect 449 -172 465 -138
rect 591 -172 607 -138
rect 641 -172 657 -138
rect 783 -172 799 -138
rect 833 -172 849 -138
rect -1091 -240 -1057 -178
rect 1057 -240 1091 -178
rect -1091 -274 -995 -240
rect 995 -274 1091 -240
<< viali >>
rect -833 138 -799 172
rect -641 138 -607 172
rect -449 138 -415 172
rect -257 138 -223 172
rect -65 138 -31 172
rect 127 138 161 172
rect 319 138 353 172
rect 511 138 545 172
rect 703 138 737 172
rect 895 138 929 172
rect -977 -88 -943 88
rect -881 -88 -847 88
rect -785 -88 -751 88
rect -689 -88 -655 88
rect -593 -88 -559 88
rect -497 -88 -463 88
rect -401 -88 -367 88
rect -305 -88 -271 88
rect -209 -88 -175 88
rect -113 -88 -79 88
rect -17 -88 17 88
rect 79 -88 113 88
rect 175 -88 209 88
rect 271 -88 305 88
rect 367 -88 401 88
rect 463 -88 497 88
rect 559 -88 593 88
rect 655 -88 689 88
rect 751 -88 785 88
rect 847 -88 881 88
rect 943 -88 977 88
rect -929 -172 -895 -138
rect -737 -172 -703 -138
rect -545 -172 -511 -138
rect -353 -172 -319 -138
rect -161 -172 -127 -138
rect 31 -172 65 -138
rect 223 -172 257 -138
rect 415 -172 449 -138
rect 607 -172 641 -138
rect 799 -172 833 -138
<< metal1 >>
rect -845 172 -787 178
rect -845 138 -833 172
rect -799 138 -787 172
rect -845 132 -787 138
rect -653 172 -595 178
rect -653 138 -641 172
rect -607 138 -595 172
rect -653 132 -595 138
rect -461 172 -403 178
rect -461 138 -449 172
rect -415 138 -403 172
rect -461 132 -403 138
rect -269 172 -211 178
rect -269 138 -257 172
rect -223 138 -211 172
rect -269 132 -211 138
rect -77 172 -19 178
rect -77 138 -65 172
rect -31 138 -19 172
rect -77 132 -19 138
rect 115 172 173 178
rect 115 138 127 172
rect 161 138 173 172
rect 115 132 173 138
rect 307 172 365 178
rect 307 138 319 172
rect 353 138 365 172
rect 307 132 365 138
rect 499 172 557 178
rect 499 138 511 172
rect 545 138 557 172
rect 499 132 557 138
rect 691 172 749 178
rect 691 138 703 172
rect 737 138 749 172
rect 691 132 749 138
rect 883 172 941 178
rect 883 138 895 172
rect 929 138 941 172
rect 883 132 941 138
rect -983 88 -937 100
rect -983 -88 -977 88
rect -943 -88 -937 88
rect -983 -100 -937 -88
rect -887 88 -841 100
rect -887 -88 -881 88
rect -847 -88 -841 88
rect -887 -100 -841 -88
rect -791 88 -745 100
rect -791 -88 -785 88
rect -751 -88 -745 88
rect -791 -100 -745 -88
rect -695 88 -649 100
rect -695 -88 -689 88
rect -655 -88 -649 88
rect -695 -100 -649 -88
rect -599 88 -553 100
rect -599 -88 -593 88
rect -559 -88 -553 88
rect -599 -100 -553 -88
rect -503 88 -457 100
rect -503 -88 -497 88
rect -463 -88 -457 88
rect -503 -100 -457 -88
rect -407 88 -361 100
rect -407 -88 -401 88
rect -367 -88 -361 88
rect -407 -100 -361 -88
rect -311 88 -265 100
rect -311 -88 -305 88
rect -271 -88 -265 88
rect -311 -100 -265 -88
rect -215 88 -169 100
rect -215 -88 -209 88
rect -175 -88 -169 88
rect -215 -100 -169 -88
rect -119 88 -73 100
rect -119 -88 -113 88
rect -79 -88 -73 88
rect -119 -100 -73 -88
rect -23 88 23 100
rect -23 -88 -17 88
rect 17 -88 23 88
rect -23 -100 23 -88
rect 73 88 119 100
rect 73 -88 79 88
rect 113 -88 119 88
rect 73 -100 119 -88
rect 169 88 215 100
rect 169 -88 175 88
rect 209 -88 215 88
rect 169 -100 215 -88
rect 265 88 311 100
rect 265 -88 271 88
rect 305 -88 311 88
rect 265 -100 311 -88
rect 361 88 407 100
rect 361 -88 367 88
rect 401 -88 407 88
rect 361 -100 407 -88
rect 457 88 503 100
rect 457 -88 463 88
rect 497 -88 503 88
rect 457 -100 503 -88
rect 553 88 599 100
rect 553 -88 559 88
rect 593 -88 599 88
rect 553 -100 599 -88
rect 649 88 695 100
rect 649 -88 655 88
rect 689 -88 695 88
rect 649 -100 695 -88
rect 745 88 791 100
rect 745 -88 751 88
rect 785 -88 791 88
rect 745 -100 791 -88
rect 841 88 887 100
rect 841 -88 847 88
rect 881 -88 887 88
rect 841 -100 887 -88
rect 937 88 983 100
rect 937 -88 943 88
rect 977 -88 983 88
rect 937 -100 983 -88
rect -941 -138 -883 -132
rect -941 -172 -929 -138
rect -895 -172 -883 -138
rect -941 -178 -883 -172
rect -749 -138 -691 -132
rect -749 -172 -737 -138
rect -703 -172 -691 -138
rect -749 -178 -691 -172
rect -557 -138 -499 -132
rect -557 -172 -545 -138
rect -511 -172 -499 -138
rect -557 -178 -499 -172
rect -365 -138 -307 -132
rect -365 -172 -353 -138
rect -319 -172 -307 -138
rect -365 -178 -307 -172
rect -173 -138 -115 -132
rect -173 -172 -161 -138
rect -127 -172 -115 -138
rect -173 -178 -115 -172
rect 19 -138 77 -132
rect 19 -172 31 -138
rect 65 -172 77 -138
rect 19 -178 77 -172
rect 211 -138 269 -132
rect 211 -172 223 -138
rect 257 -172 269 -138
rect 211 -178 269 -172
rect 403 -138 461 -132
rect 403 -172 415 -138
rect 449 -172 461 -138
rect 403 -178 461 -172
rect 595 -138 653 -132
rect 595 -172 607 -138
rect 641 -172 653 -138
rect 595 -178 653 -172
rect 787 -138 845 -132
rect 787 -172 799 -138
rect 833 -172 845 -138
rect 787 -178 845 -172
<< properties >>
string FIXED_BBOX -1074 -257 1074 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.15 m 1 nf 20 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
